(** This module reexports all the modules in Logic.Effects.*. *)

From Metaprog.Logic.Effects Require Export Print Fail Iter Rec Evar.
