(** This module re-exports all effects. *)

From Metaprog.Control.Effects Require Export Print Fail Iter Rec Evar.