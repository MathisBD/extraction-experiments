(** This module loads the ocaml plugin. *)

Declare ML Module "extraction-experiments.plugin".