(** This module loads the OCaml plugin against which the extracted code is linked. *)

Declare ML Module "extraction-experiments.plugin".
